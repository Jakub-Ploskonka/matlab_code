Roznicowy

*model scalonego tranzystora bipolarnego
.MODEL trNPN NPN BF=80 BR=1 IS=1.0E-14 RB=100 VA=50 TF=0.3N TR=6.0N
+ CCS=2.0P CJE=3.0P CJC=2.0P KF=6.6E-16 AF=1
*

vcc vcc 0 5
vee vee 0 -5

q1 vcc we1 e trnpn
q2 vcc we2 e trnpn
q3 e b34 vee trnpn
q4 b34 b34 vee trnpn

iee vcc b34 0.5m

vwe1 we1 0 {cm+diff}
vwe2 we2 0 {cm-diff}

.param cm=0
.param diff=0

.dc param vcc -1 1 1m
.dc param diff -100m 100m 1m
.probe
.end